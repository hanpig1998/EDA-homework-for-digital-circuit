library verilog;
use verilog.vl_types.all;
entity mul2_vlg_vec_tst is
end mul2_vlg_vec_tst;
